module TopLevel #(parameter N = 32)(input logic clk,
												output logic [31:0]z_RD1,
												output logic [31:0]z_RD2,
												output logic [12:0]z_MD,
												output logic [31:0]z_ALU_out,
												output logic [31:0]z_ALU_in1,
												output logic [31:0]z_ALU_in2,
												output logic [31:0]z_RF_WD);
												
												
	
	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	//////////////////////////////////////////////////////////////ALU///////////////////////////////////////////////////////////////	
	logic ALU_cmp_out;
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	///////////////////////////////////////////////Multiplexor Before ALU input IN2/////////////////////////////////////////////////	
	logic [31:0]ALU_IN2_in;
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	///////////////////////////////////////////////////////Register File////////////////////////////////////////////////////////////	
	logic [31:0]RF_RD1_out;
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	//////////////////////////////////////////Multiplexor Before Register File input WD/////////////////////////////////////////////	
	logic [31:0]LDIT_out;
	logic [31:0]RAM_out;
	logic [31:0]ALU_out;
	logic [31:0]RF_RD2_out;
	logic [31:0]RF_WD_in;
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	///////////////////////////////////////////////////////MAIN DECODER/////////////////////////////////////////////////////////////	
	logic [12:0]state;
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	///////////////////////////////////////////////////////ROM//////////////////////////////////////////////////////////////////////	
	logic [10:0]ROM_in;
	logic [31:0]ROM_out;
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	logic reset;
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	Reset res(.clk(clk),.reset(reset));
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	ROM rom_instance(.adr(ROM_in), .dout(ROM_out));
	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	MainDecoder mainDecoder_instance(.cmd(ROM_out[4:0]), .out(state));
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	decoderLDI decLDI(.data(ROM_out[31:16]), .switch(state[7]), .dataOut(LDIT_out));
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	RegisterFile registerFile_instance(.clk(clk), .reset(reset), .WE(state[1]), .A1(ROM_out[9:5]), .A2(ROM_out[14:10]),
										.WD(RF_WD_in), .RD1(RF_RD1_out), .RD2(RF_RD2_out));
	
	always_comb begin
		case(state[3:2])
			2'b11:	RF_WD_in = RF_RD2_out;
			2'b10:	RF_WD_in = ALU_out;
			2'b01:	RF_WD_in = RAM_out;
			2'b00:	RF_WD_in = LDIT_out;
		endcase
	end	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	RAM ram_instance(.clk(clk), .we(state[0]), .addr(RF_RD2_out[7:0]), .dataIn(RF_RD1_out), .dataOut(RAM_out));
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	always_comb begin
		case(state[6:5])
			2'b11:	ALU_IN2_in = 32'd0;
			2'b10:	ALU_IN2_in = {27'd0,ROM_out[14:10]};
			2'b01:	ALU_IN2_in = RF_RD2_out;
			2'b00:	ALU_IN2_in = 32'd0;
		endcase
	end
	ALU alu_instance(.dataIn0(RF_RD1_out), .dataIn1(ALU_IN2_in), .ctrlALU(state[11:8]), .cmp(ALU_cmp_out), .dataOut(ALU_out));
	
	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	InstructionCounter IC(.clk(clk), .reset(reset), .shift(ROM_out[31:16]), .MD_mux0_ctrl(state[4]), 
									.MD_mux1_ctrl(state[12]), .ALU_mux1_ctrl(ALU_cmp_out), .out(ROM_in));
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	assign ROM_out[15] = 1'd0;
	always_comb begin
		z_RD1 <= RF_RD1_out;
		z_RD2 <= RF_RD2_out;
		z_MD <= state;
		z_ALU_out <= ALU_out;
		z_ALU_in1 <= RF_RD1_out;
		z_ALU_in2 <= ALU_IN2_in;
		z_RF_WD <= RF_WD_in;
	end

endmodule 















